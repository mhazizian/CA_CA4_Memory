// LENGHTs

`define ADDRESS_LEN 		15
`define TAG_LEN				1
`define WORD_LEN			32
`define CACHE_INDEX_LEN		12

`define CACHE_BLOCK_LEN		130
`define CACHE_CAPACITY		4096
`define MEM_CAPACITY		32768
